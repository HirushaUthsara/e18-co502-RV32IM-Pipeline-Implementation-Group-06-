
`timescale 1ns/100ps

module BRANCH_HAZZARDS(ID_PC, ALU_PC, RESET, ID_BRANCH, ALU_BRANCH, ALU_BRANCH_RESULT, FLUSH, EARLY_PREDICT, TAKE_BRANCH);

    input [2:0] ID_PC, ALU_PC;
    input RESET, ID_BRANCH, ALU_BRANCH, ALU_BRANCH_RESULT;
    output reg FLUSH, EARLY_PREDICT, TAKE_BRANCH;

    reg [1:0] PREDICTION[0:7];

    parameter BRANCH_TAKEN_STRONG = 2'b00, BRANCH_TAKEN_WEAK = 2'b01, BRANCH_NOTTAKEN_WEAK = 2'b10, BRANCH_NOTTAKEN_STRONG = 2'b11;

    // Logic for ALU_BRANCH prediction
    always @(*) begin
        if (ALU_BRANCH) begin
            case (PREDICTION[ALU_PC])
                BRANCH_TAKEN_STRONG:
                    if (ALU_BRANCH_RESULT) begin
                        PREDICTION[ALU_PC] = 2'b00;
                        FLUSH = 1'b0;
                    end
                    else begin
                        PREDICTION[ALU_PC] = 2'b01;
                        FLUSH = 1'b1;
                        EARLY_PREDICT = 1'b1;
                    end
                BRANCH_TAKEN_WEAK:
                    if (ALU_BRANCH_RESULT) begin
                        PREDICTION[ALU_PC] = 2'b00;
                        FLUSH = 1'b0;
                    end
                    else begin
                        PREDICTION[ALU_PC] = 2'b10;
                        FLUSH = 1'b1;
                        EARLY_PREDICT = 1'b1;
                    end
                BRANCH_NOTTAKEN_WEAK:
                    if (ALU_BRANCH_RESULT) begin
                        PREDICTION[ALU_PC] = 2'b01;
                        FLUSH = 1'b1;
                        EARLY_PREDICT = 1'b0;
                    end
                    else begin
                        PREDICTION[ALU_PC] = 2'b11;
                        FLUSH = 1'b0;
                    end
                BRANCH_NOTTAKEN_STRONG:
                    if (ALU_BRANCH_RESULT) begin
                        PREDICTION[ALU_PC] = 2'b10;
                        FLUSH = 1'b1;
                        EARLY_PREDICT = 1'b0;
                    end
                    else begin
                        PREDICTION[ALU_PC] = 2'b11;
                        FLUSH = 1'b0;
                    end
            endcase
        end
        else begin
            FLUSH = 1'b0;
        end
    end

    // Logic for ID_BRANCH prediction
    always @(*) begin
        if (ID_BRANCH) begin
            case (PREDICTION[ID_PC])
                BRANCH_TAKEN_STRONG:
                    TAKE_BRANCH = 1'b1;
                BRANCH_TAKEN_WEAK:
                    TAKE_BRANCH = 1'b1;
                BRANCH_NOTTAKEN_WEAK:
                    TAKE_BRANCH = 1'b0;
                BRANCH_NOTTAKEN_STRONG:
                    TAKE_BRANCH = 1'b0;
            endcase
        end
        else begin
            TAKE_BRANCH = 1'b0;
        end
    end

    // Initializing all branch decisions to BRANCH_TAKEN_STRONG state
    integer i;
    always @(RESET) begin
        FLUSH = 1'b0;
        for (i = 0; i < 8; i = i + 1) begin
            PREDICTION[i] = 2'b00;
        end
    end

endmodule


/*
ID_PC: The program counter (PC) value at the Instruction Decode (ID) stage. It represents the address of the current instruction being processed in the pipeline.

ALU_PC: The program counter (PC) value at the Arithmetic Logic Unit (ALU) stage. It represents the address of the instruction being processed by the ALU.

RESET: A control signal that initiates a reset operation in the pipeline. When RESET is asserted, the pipeline stages are cleared, and the pipeline is brought to an initial state.

ID_STAGE_BRANCH: A control signal indicating whether a branch instruction is encountered in the Instruction Decode (ID) stage. It is typically generated by the instruction decoder based on the opcode and determines if the current instruction is a branch instruction.

ALU_STAGE_BRANCH: A control signal indicating whether a branch instruction is being processed in the Arithmetic Logic Unit (ALU) stage. It is typically generated based on the type of branch instruction and determines if the current instruction is a branch instruction being executed by the ALU.

ALU_STAGE_BRANCH_RESULT: A signal that holds the result of the branch operation performed by the ALU. It represents the outcome of the branch instruction, such as whether the branch is taken or not.

FLUSH: A control signal used to flush or discard instructions in the pipeline. When FLUSH is asserted, it indicates that the instructions currently in the pipeline should be invalidated or cleared.

EARLY_PREDICTION: A technique used in branch prediction algorithms to predict the outcome of a branch instruction before it is executed. This signal indicates whether an early prediction is made for the branch instruction.

TAKE_BRANCH: A control signal indicating whether the branch instruction should be taken. It is typically based on the branch result from the ALU and the branch prediction. When TAKE_BRANCH is asserted, it indicates that the branch should be taken and the pipeline needs to be redirected to the target address specified by the branch instruction.

This module represents a branch predictor. Here's a summary of its functionality:

Input Ports:

ID_PC and ALU_PC: Current program counters for the ID and ALU stages.
RESET: Reset signal.
ID_BRANCH and ALU_BRANCH: Branch signals indicating the presence of a branch instruction in the ID and ALU stages, respectively.
ALU_BRANCH_RESULT: Result of the branch prediction from the ALU stage.
Output Ports:

FLUSH: Signal indicating whether the pipeline needs to be flushed.
EARLY_PREDICT: Signal indicating whether early branch prediction is enabled.
TAKE_BRANCH: Signal indicating whether the branch should be taken.
Internal Signals:

PREDICTION: Array of 2-bit registers representing the prediction state for different program counters.
BRANCH_TAKEN_STRONG, BRANCH_TAKEN_WEAK, BRANCH_NOTTAKEN_WEAK, BRANCH_NOTTAKEN_STRONG: Parameter values representing different branch prediction states.
Functionality:

The module uses two separate always blocks to handle the branch prediction for the ALU stage and ID stage.
In the ALU stage branch prediction, the module checks the current prediction state stored in PREDICTION[ALU_PC] and evaluates the branch result (ALU_BRANCH_RESULT).
Depending on the prediction state and branch result, the module updates the prediction state, sets the FLUSH signal accordingly, and determines the EARLY_PREDICT value.
Similarly, in the ID stage branch prediction, the module checks the current prediction state stored in PREDICTION[ID_PC] and sets the TAKE_BRANCH signal based on the prediction state.
The RESET signal is used to initialize all branch predictions to the BRANCH_TAKEN_STRONG state in the always @(RESET) block.
Overall, this module implements a branch predictor that uses prediction states and branch results to determine whether to take the branch and whether to flush the pipeline.
*/