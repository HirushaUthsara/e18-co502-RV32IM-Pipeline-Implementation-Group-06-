`timescale  1ns/100ps

`include "../Adder/Adder.v"
`include "../ALU/ALU.v"
`include "../Branch_Jump/Branch_Jump.v"
`include "../Control_unit/ControlUnit.v"
`include "../Data_Memory/Data_Memory.v"
`include "../Data_Memory/Data_Correcting.v"
`include "../DataCache/data_cache.v"
//`include "../ImmediateGenerator/ImmediateGenarator.v"
//`include "../Instruction_fetch_module/InstructionFetch.v"
`include "../InstructionCache/instruction_cache.v"
`include "../InstructionMemory/InstructionMemory.v"
`include "../Mux/MUX.v"
`include "../PC/PC.v"
`include "../Pipeline_Registers/Pipeline_Registers.v"
`include "../Register_File/RegisterFile.v"
`include "../Sign_Zero_Extend/Sign_Zero_Extend.v"



module CPU(CLK, RESET);

// port declaration
input RESET, CLK; 

wire WRITE_REG, MUXPC_SELECT, MUXIMM_SELECT, MUXJAL_SELECT, MUXDATAMEM_SELECT, WRITE_ENABLE, MEM_READ, MEM_WRITE, BRANCH, JUMP;
wire [31:0] INSTRUCTION, IN_REG, OUT1_REG, OUT2_REG, SIGN_ZERO_EXTEND,  PC_DIRECT_OUT_IN, PC_PLUS_4_OUT_IN;
wire [4:0] MEM_WB_INADDRESS, ALUOP;
wire[2:0] MUXIMMTYPE_SELECT;

// ID/EX and EX/MEM stage wires
wire EQ_FLAG, LT_FLAG, LTU_FLAG, PC_MUX_CONTROL, REG_FLUSH;
wire [31:0] DATA1, DATA2, RESULT_ALU, MUXJAL_OUT, BRANCH_OR_JUMP_ADDR;

// EX/MEM and MEM/WB stage wires
wire MEM_BUSYWAIT, MEM_MEM_READ, MEM_MEM_WRITE; 
wire [27:0] MEM_BLOCK_ADDR;
wire [31:0] CACHE_READ_OUT;
wire [127:0] DATA_MEM_READ_OUT, DATA_MEM_WRITE_OUT;

// MEM/WB and IF/ID stage
wire [31:0] PC, PC_PLUS_4, PC_MUX_OUT;


// ID_EX Register Outputs
wire WRITE_ENABLE_OUT, MUXDATAMEM_SELECT_OUT, MEM_READ_OUT, MEM_WRITE_OUT, MUXJAL_SELECT_OUT, MUXIMM_SELECT_OUT, MUXPC_SELECT_OUT, BRANCH_OUT, JUMP_OUT;
wire [2:0] FUNCT3_OUT;
wire [4:0] ALUOP_OUT, RD_OUT;
wire [31:0] PC_DIRECT_OUT_OUT, SIGN_ZERO_EXTEND_OUT, PC_PLUS_4_OUT_OUT, OUT1_OUT, OUT2_OUT;

// EX_MEM Register Outputs
wire WRITE_ENABLE_OUT_EX_MEM,  MUXDATAMEM_SELECT_OUT_EX_MEM, MEM_READ_OUT_EX_MEM, MEM_WRITE_OUT_EX_MEM;
wire [2:0] FUNCT3_OUT_EX_MEM;
wire [4:0] RD_OUT_EX_MEM;
wire [31:0] MUXJAL_OUT_EX_MEM, OUT2_OUT_EX_MEM;

// MEM_WB Register Outputs
wire  MUXDATAMEM_SELECT_OUT_MEM_WB;
wire [31:0] CACHE_READ_OUT_MEM_WB, MUXJAL_OUT_MEM_WB, DATA_CORRECTING_OUT, TO_DATA_MEM;

wire [31:0] READINST;
wire [27:0] MEM_ADDRESS_TO_CACHE;
wire [127:0] MEM_READINST;
wire I_BUSYWAIT, I_MEM_READ, I_MEM_BUSYWAIT;

wire BUSYWAIT, D_BUSYWAIT;

assign BUSYWAIT = D_BUSYWAIT || I_BUSYWAIT;

// Stage 2
    register_file  regfile(MEM_WB_INADDRESS, IN_REG, INSTRUCTION[19:15], INSTRUCTION[24:20],  OUT1_REG, OUT2_REG,  WRITE_REG, CLK, RESET);
    CONTROL_UNIT controlunit(INSTRUCTION, ALUOP,  MUXIMMTYPE_SELECT, MUXPC_SELECT, MUXIMM_SELECT, MUXJAL_SELECT, MUXDATAMEM_SELECT, WRITE_ENABLE, MEM_READ, MEM_WRITE, BRANCH, JUMP);
    Sign_Zero_Extend signZeroExtend(INSTRUCTION,MUXIMMTYPE_SELECT, SIGN_ZERO_EXTEND );
    PIPEREG2 reg2(CLK,REG_FLUSH,WRITE_ENABLE,MUXDATAMEM_SELECT,
    MEM_READ,MEM_WRITE,MUXJAL_SELECT,ALUOP,MUXIMM_SELECT,
    MUXPC_SELECT,BRANCH,JUMP,PC_DIRECT_OUT_IN,SIGN_ZERO_EXTEND,
    PC_PLUS_4_OUT_IN,OUT1_REG,OUT2_REG, INSTRUCTION[11:7],INSTRUCTION[14:12],
    WRITE_ENABLE_OUT,MUXDATAMEM_SELECT_OUT,MEM_READ_OUT,MEM_WRITE_OUT,
    MUXJAL_SELECT_OUT,ALUOP_OUT,MUXIMM_SELECT_OUT,MUXPC_SELECT_OUT,BRANCH_OUT,
    JUMP_OUT,PC_DIRECT_OUT_OUT,SIGN_ZERO_EXTEND_OUT,PC_PLUS_4_OUT_OUT,OUT1_OUT,
    OUT2_OUT,RD_OUT,FUNCT3_OUT,BUSYWAIT);

// stage 3
    MUX_A Mux1(OUT1_OUT, PC_DIRECT_OUT_OUT, DATA1, MUXPC_SELECT_OUT);
    MUX_A Mux2(OUT2_OUT, SIGN_ZERO_EXTEND_OUT, DATA2, MUXIMM_SELECT_OUT);
    ALU alu(DATA1, DATA2, RESULT_ALU, ALUOP_OUT, EQ_FLAG, LT_FLAG, LTU_FLAG);
    MUX_A Mux3(RESULT_ALU, PC_PLUS_4_OUT_OUT, MUXJAL_OUT, MUXJAL_SELECT_OUT);
    BRANCH_JUMP branchjump(RESET,RESULT_ALU, SIGN_ZERO_EXTEND_OUT, FUNCT3_OUT, BRANCH_OUT, JUMP_OUT, EQ_FLAG, LT_FLAG, LTU_FLAG, BRANCH_OR_JUMP_ADDR, PC_MUX_CONTROL, REG_FLUSH);
    PIPEREG3 reg3(CLK, REG_FLUSH, WRITE_ENABLE_OUT, MUXDATAMEM_SELECT_OUT, MEM_READ_OUT,
    MEM_WRITE_OUT, MUXJAL_OUT, OUT2_OUT, RD_OUT, FUNCT3_OUT, 
    WRITE_ENABLE_OUT_EX_MEM,  MUXDATAMEM_SELECT_OUT_EX_MEM, MEM_READ_OUT_EX_MEM, 
    MEM_WRITE_OUT_EX_MEM, MUXJAL_OUT_EX_MEM, OUT2_OUT_EX_MEM, RD_OUT_EX_MEM, 
    FUNCT3_OUT_EX_MEM, BUSYWAIT);


// stage 4
    DATA_CACHE datacache(CLK, RESET, MEM_READ_OUT_EX_MEM, MEM_WRITE_OUT_EX_MEM, MUXJAL_OUT_EX_MEM, TO_DATA_MEM, 
    MEM_BUSYWAIT, DATA_MEM_READ_OUT, CACHE_READ_OUT, MEM_MEM_READ, MEM_MEM_WRITE, D_BUSYWAIT, MEM_BLOCK_ADDR, DATA_MEM_WRITE_OUT);
    DATA_MEMORY dmem(CLK, RESET, MEM_MEM_READ, MEM_MEM_WRITE, MEM_BLOCK_ADDR, DATA_MEM_WRITE_OUT, DATA_MEM_READ_OUT, MEM_BUSYWAIT);
    DATA_CORRECTING datacorrecting(FUNCT3_OUT_EX_MEM, CACHE_READ_OUT,DATA_CORRECTING_OUT, TO_DATA_MEM, OUT2_OUT_EX_MEM);
    PIPEREG4 reg4(CLK, REG_FLUSH, WRITE_ENABLE_OUT_EX_MEM,  MUXDATAMEM_SELECT_OUT_EX_MEM, DATA_CORRECTING_OUT, 
    MUXJAL_OUT_EX_MEM, RD_OUT_EX_MEM, WRITE_REG, MUXDATAMEM_SELECT_OUT_MEM_WB, 
    CACHE_READ_OUT_MEM_WB, MUXJAL_OUT_MEM_WB, MEM_WB_INADDRESS, BUSYWAIT);

// stage 5-1
    MUX_A Mux4(MUXJAL_OUT_MEM_WB, CACHE_READ_OUT_MEM_WB, IN_REG, MUXDATAMEM_SELECT_OUT_EX_MEM);
    MUX_A Mux(PC_PLUS_4, BRANCH_OR_JUMP_ADDR, PC_MUX_OUT, PC_MUX_CONTROL);
    PC pc(PC_MUX_OUT, PC, RESET, CLK, BUSYWAIT);
    adder_4 pcadder(PC, PC_PLUS_4);
    instruction_cache instructioncache(CLK,RESET, PC, READINST,   I_BUSYWAIT, MEM_ADDRESS_TO_CACHE, I_MEM_READ, MEM_READINST, I_MEM_BUSYWAIT);
    INSTRUCTION_MEMORY instmem( CLK,I_MEM_READ,MEM_ADDRESS_TO_CACHE,MEM_READINST,I_MEM_BUSYWAIT);
    PIPEREG1 reg1(CLK,REG_FLUSH,READINST,PC_PLUS_4,PC,INSTRUCTION,PC_PLUS_4_OUT_IN,PC_DIRECT_OUT_IN,BUSYWAIT);

endmodule


module cpu_tb;

    reg CLK, RESET;

    CPU cpu(CLK, RESET);
	
    initial
    begin
    
        // generate files needed to plot the waveform using GTKWave
        $dumpfile("cpu_wavedata.vcd");
	    $dumpvars(0, cpu_tb);
        
        CLK = 1'b0;
		RESET = 1'b0;
		RESET = 1'b1;
		#4;
		RESET = 1'b0;
		
		#15000;
		$finish;
        
    end
    

// clock genaration.
always begin
    #3 CLK = ~CLK;
end

endmodule